module InstrDecoder(output reg [2:0] o_ImmSrc,
                    input      [6:0] i_Op);

//`include "src/IType.v"
localparam [2:0] NO = 3'd0,
                 RT = 3'd1,
                 IT = 3'd2,
                 ST = 3'd3,
                 BT = 3'd4,
                 UT = 3'd5,
                 JT = 3'd6;

always @(*)
begin
	casez (i_Op)
		7'b011_0011: o_ImmSrc = RT;

		7'b001_0011: o_ImmSrc = IT;
		7'b000_0011: o_ImmSrc = IT;
		7'b110_0111: o_ImmSrc = IT;
		7'b111_0011: o_ImmSrc = IT;

		7'b010_0011: o_ImmSrc = ST;
		7'b110_0011: o_ImmSrc = BT;
		7'b110_1111: o_ImmSrc = JT;
		7'b0?1_0111: o_ImmSrc = UT;
		default:     o_ImmSrc = NO;
	endcase
end

endmodule

