module IssueQueue(output [] o_issue);




endmodule

